magic
tech scmos
timestamp 1669664801
<< metal1 >>
rect -1691 836 -1631 840
rect -1719 829 -1631 833
rect -1719 377 -1715 829
rect -1565 826 1586 830
rect -781 736 584 737
rect -781 733 1586 736
rect 544 732 1586 733
rect -1691 380 -1631 384
rect -781 382 -636 386
rect -1719 373 -1631 377
rect -1719 291 -1715 373
rect -1565 370 -1492 374
rect -1690 294 -1630 298
rect -1719 287 -1631 291
rect -1719 205 -1715 287
rect -1565 284 -1514 288
rect -1498 287 -1492 370
rect -1519 274 -1514 284
rect -1519 264 -1492 274
rect -1515 222 -1492 232
rect -1691 208 -1631 212
rect -1719 201 -1631 205
rect -1515 202 -1510 222
rect -1719 152 -1715 201
rect -1565 198 -1510 202
rect -1499 156 -1492 209
rect -781 4 -698 8
rect -1686 -93 -1626 -89
rect -1715 -100 -1626 -96
rect -1715 -182 -1711 -100
rect -1560 -103 -1497 -99
rect -1504 -162 -1497 -103
rect -1504 -170 -1491 -162
rect -1686 -179 -1626 -175
rect -1715 -186 -1626 -182
rect -1715 -268 -1711 -186
rect -1560 -189 -1501 -185
rect -1506 -196 -1501 -189
rect -1506 -204 -1491 -196
rect -1517 -233 -1491 -225
rect -1686 -265 -1626 -261
rect -1715 -272 -1626 -268
rect -1517 -271 -1511 -233
rect -1715 -354 -1711 -272
rect -1560 -275 -1511 -271
rect -1500 -271 -1491 -263
rect -1686 -351 -1626 -347
rect -1715 -358 -1626 -354
rect -1500 -357 -1494 -271
rect -1715 -390 -1711 -358
rect -1560 -361 -1494 -357
rect -781 -371 -745 -367
rect -755 -627 -745 -371
rect -707 -585 -698 4
rect -646 -562 -636 382
rect 325 -126 1586 -122
rect 1573 -127 1586 -126
rect 325 -477 457 -473
rect -646 -572 -386 -562
rect -707 -595 -386 -585
rect -756 -638 -385 -627
rect -781 -648 -773 -641
rect -780 -650 -773 -648
rect -780 -660 -386 -650
rect 325 -855 395 -851
rect -580 -952 -520 -948
rect -609 -959 -520 -955
rect -609 -1041 -605 -959
rect -454 -962 -391 -958
rect -398 -1021 -391 -962
rect -398 -1029 -385 -1021
rect -580 -1038 -520 -1034
rect -609 -1045 -520 -1041
rect -609 -1127 -605 -1045
rect -454 -1048 -395 -1044
rect -400 -1055 -395 -1048
rect -400 -1063 -385 -1055
rect -411 -1092 -385 -1084
rect -580 -1124 -520 -1120
rect -609 -1131 -520 -1127
rect -411 -1130 -405 -1092
rect -609 -1213 -605 -1131
rect -454 -1134 -405 -1130
rect -394 -1130 -385 -1122
rect -580 -1210 -520 -1206
rect -609 -1217 -520 -1213
rect -394 -1216 -388 -1130
rect -609 -1249 -605 -1217
rect -454 -1220 -388 -1216
rect 325 -1230 348 -1226
rect 338 -1486 348 -1230
rect 386 -1444 395 -855
rect 447 -1421 457 -477
rect 1418 -985 1586 -981
rect 1418 -1336 1586 -1332
rect 447 -1431 707 -1421
rect 386 -1454 707 -1444
rect 337 -1497 708 -1486
rect 325 -1509 329 -1499
rect 325 -1519 707 -1509
rect 1418 -1714 1586 -1710
rect 513 -1811 573 -1807
rect 484 -1818 573 -1814
rect 484 -1900 488 -1818
rect 639 -1821 702 -1817
rect 695 -1880 702 -1821
rect 695 -1888 708 -1880
rect 513 -1897 573 -1893
rect 484 -1904 573 -1900
rect 484 -1986 488 -1904
rect 639 -1907 698 -1903
rect 693 -1914 698 -1907
rect 693 -1922 708 -1914
rect 682 -1951 708 -1943
rect 513 -1983 573 -1979
rect 484 -1990 573 -1986
rect 682 -1989 688 -1951
rect 484 -2072 488 -1990
rect 639 -1993 688 -1989
rect 699 -1989 708 -1981
rect 513 -2069 573 -2065
rect 484 -2076 573 -2072
rect 699 -2075 705 -1989
rect 484 -2108 488 -2076
rect 639 -2079 705 -2075
rect 1418 -2089 1586 -2085
rect 1418 -2367 1586 -2358
use AND  AND_11
timestamp 1669664801
transform 1 0 573 0 1 -2106
box 0 0 66 83
use AND  AND_14
timestamp 1669664801
transform 1 0 573 0 1 -1848
box 0 0 66 83
use AND  AND_13
timestamp 1669664801
transform 1 0 573 0 1 -1934
box 0 0 66 83
use AND  AND_12
timestamp 1669664801
transform 1 0 573 0 1 -2020
box 0 0 66 83
use AND  AND_9
timestamp 1669664801
transform 1 0 -520 0 1 -1247
box 0 0 66 83
use AND  AND_10
timestamp 1669664801
transform 1 0 -520 0 1 -1161
box 0 0 66 83
use AND  AND_8
timestamp 1669664801
transform 1 0 -520 0 1 -1075
box 0 0 66 83
use AND  AND_3
timestamp 1669664801
transform 1 0 -520 0 1 -989
box 0 0 66 83
use AND  AND_4
timestamp 1669664801
transform 1 0 -1626 0 1 -302
box 0 0 66 83
use AND  AND_5
timestamp 1669664801
transform 1 0 -1626 0 1 -388
box 0 0 66 83
use AND  AND_6
timestamp 1669664801
transform 1 0 -1626 0 1 -216
box 0 0 66 83
use AND  AND_7
timestamp 1669664801
transform 1 0 -1626 0 1 -130
box 0 0 66 83
use AND  AND_2
timestamp 1669664801
transform 1 0 -1631 0 1 171
box 0 0 66 83
use AND  AND_1
timestamp 1669664801
transform 1 0 -1631 0 1 257
box 0 0 66 83
use AND  AND_0
timestamp 1669664801
transform 1 0 -1631 0 1 343
box 0 0 66 83
use Adder_4  Adder_4_0
timestamp 1668116499
transform 0 -1 -874 1 0 -266
box -382 -93 1069 618
use Adder_4  Adder_4_1
timestamp 1668116499
transform 0 -1 232 1 0 -1125
box -382 -93 1069 618
use AND  AND_15
timestamp 1669664801
transform 1 0 -1631 0 1 799
box 0 0 66 83
use Adder_4  Adder_4_2
timestamp 1668116499
transform 0 -1 1325 1 0 -1984
box -382 -93 1069 618
<< labels >>
rlabel metal1 1580 826 1580 830 7 P0
rlabel metal1 1581 732 1581 736 7 P1
rlabel metal1 1580 -127 1580 -123 7 P2
rlabel metal1 1581 -985 1581 -981 7 P3
rlabel metal1 1581 -1336 1581 -1332 7 P4
rlabel metal1 1579 -1714 1579 -1710 7 P5
rlabel metal1 1581 -2089 1581 -2085 7 P6
rlabel metal1 1573 -2366 1580 -2365 1 P7
rlabel metal1 -1494 162 -1493 180 7 gnd
rlabel metal1 -1679 208 -1678 212 7 B3
rlabel metal1 -1677 294 -1676 298 7 B2
rlabel metal1 -1680 380 -1679 384 7 B1
rlabel metal1 -1675 836 -1674 840 7 B0
rlabel metal1 -1717 157 -1716 166 3 A0
rlabel metal1 -1668 -351 -1668 -347 7 B3
rlabel metal1 -1670 -265 -1670 -261 7 B2
rlabel metal1 -1672 -179 -1672 -175 7 B1
rlabel metal1 -1671 -93 -1671 -89 7 B0
rlabel metal1 -558 -1210 -558 -1206 7 B3
rlabel metal1 -559 -1124 -559 -1120 7 B2
rlabel metal1 -560 -1038 -560 -1034 7 B1
rlabel metal1 -561 -952 -561 -948 7 B0
rlabel metal1 531 -2069 531 -2065 7 B3
rlabel metal1 530 -1983 530 -1979 7 B2
rlabel metal1 528 -1897 528 -1893 7 B1
rlabel metal1 529 -1811 529 -1807 7 B0
rlabel metal1 486 -2100 486 -2096 7 A3
rlabel metal1 -607 -1244 -607 -1240 7 A2
rlabel metal1 -1713 -386 -1713 -382 7 A1
<< end >>
